
module test();
	wire [3:0] a = 4'hFF;
	initial begin
		$display("%d",a);
		//assign a = '1;
		//$display("%d",a);
	end

endmodule
